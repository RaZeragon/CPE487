-- Author: N/A
-- Date: 7/11/2017
-- Title: D Flip Flop
-- Code Version: N/A
-- Type: N/A
-- Availability: https://electronicstopper.blogspot.com/2017/07/d-flip-flop-in-vhdl-with-testbench.html

library ieee;
use ieee.std_logic_1164.all;

entity DFF is 
port( din: in std_logic;
	clk: in std_logic;
	rst: in std_logic;
	dout: out std_logic);
end DFF;

architecture behavioral of DFF is
begin
	process(rst,clk,din)
	begin
		if (rst = '1') then
			dout <= '0';
		elsif (rising_edge(clk)) then
			dout <= din;
		end if;
	end process;
end behavioral;