-- Author: N/A
-- Date: 7/11/2017
-- Title: T Flip Flop
-- Code Version: N/A
-- Type: N/A
-- Availability: https://electronicstopper.blogspot.com/2017/07/t-flip-flop-in-vhdl-with-testbench.html

library ieee;
use ieee.std_logic_1164.all;

entity TFF is
	port( din: in std_logic;
		clk: in std_logic;
		rst: in std_logic;
		dout: out std_logic);
end TFF;

architecture behavioral of TFF is
begin
	process(rst, clk, din)
	begin
		if (rst = '1') then
			dout <= '0';
		elsif (rising_edge(clk)) then
			dout <= not din;
		end if;
	end process;
end behavioral;